.title KiCad schematic
.include "C:/AE/ZXCT210/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/ZXCT210/ZXCT210.LIB"
R1 /IN- /VIN {RSNS}
XU1 /VREF 0 /VSUPPLY /VIN /IN- /CNV ZXCT210
I1 /IN- 0 DC {ILOAD} 
XU2 /OUT 0 CEU4J2X7R2A103K125AE_s
R2 /CNV /OUT {ROUT}
V1 /VIN 0 DC {VIN} 
V2 /VREF 0 DC {VREF} 
V3 /VSUPPLY 0 DC {VSUPPLY} 
.end
