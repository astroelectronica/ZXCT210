.title KiCad schematic
.include "C:/AE/ZXCT210/ZXCT210.LIB"
V3 /VSUPPLY 0 DC {VSUPPLY} 
V2 /VREF 0 DC {VREF} 
V1 /VIN 0 DC {VIN} 
R1 /IN- /VIN {RSNS}
XU1 /VREF 0 /VSUPPLY /VIN /IN- /OUT ZXCT210
I1 /IN- 0 DC {ILOAD} 
.end
